`define INFO_WID  7:0
`define INFO_NUM  0:3071  // 96*32
`define COLOR_WID 4:0
