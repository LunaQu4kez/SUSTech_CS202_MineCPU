`include "Const.svh"

module Branch_Predictor (
    input  logic             clk, rst,
    input  logic [`DATA_WID] old_PC,
    output logic [`DATA_WID] new_PC
);

endmodule