`define INFO_WID  7:0
`define VGA_ADDR  11:0  // 96*32
`define COLOR_WID 4:0
