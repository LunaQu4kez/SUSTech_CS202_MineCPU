module ALU(
    input  [31:0] src1,
                  src2,
    input  [3:0]  ALUcontrol,
    output [31:0] res,
    output        zero
);




    
endmodule