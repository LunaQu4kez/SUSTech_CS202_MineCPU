module ALU (
    input [31:0]            data1, data2,
    input [3:0]             ALUop,
    output [31:0]           res,
    output                  zero
);




    
endmodule