module CPU (

);

endmodule