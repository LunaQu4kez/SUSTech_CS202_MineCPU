module ALU_Ctrl (
    input [3:0]         inst_piece1, ALUop_in,
    output [3:0]        ALUop_out
);




    
endmodule