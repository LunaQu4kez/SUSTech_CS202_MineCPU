`include "Const.svh"

module Stage_ID (

);

endmodule