`define SEG_FREQ 200000      // 500Hz
`define SEG0 8'b1111_1100    // Display '0'
`define SEG1 8'b0110_0000    // Display '1'
`define SEG2 8'b1101_1010    // Display '2'
`define SEG3 8'b1111_0010    // Display '3'
`define SEG4 8'b0110_0110    // Display '4'
`define SEG5 8'b1011_0110    // Display '5'
`define SEG6 8'b1011_1110    // Display '6'
`define SEG7 8'b1110_0000    // Display '7'
`define SEG8 8'b1111_1110    // Display '8'
`define SEG9 8'b1111_0110    // Display '9'
`define SEGA 8'b1110_1110    // Display 'A'
`define SEGB 8'b0011_1110    // Display 'B'
`define SEGC 8'b1001_1100    // Display 'C'
`define SEGD 8'b0111_1010    // Display 'D'
`define SEGE 8'b1001_1110    // Display 'E'
`define SEGF 8'b1000_1110    // Display 'F'

`define IN0 8'b00000000      // Encode of '0'
`define IN1 8'b00000001      // Encode of '1'
`define IN2 8'b00000010      // Encode of '2'
`define IN3 8'b00000011      // Encode of '3'
`define IN4 8'b00000100      // Encode of '4'
`define IN5 8'b00000101      // Encode of '5'
`define IN6 8'b00000110      // Encode of '6'
`define IN7 8'b00000111      // Encode of '7'
`define IN8 8'b00001000      // Encode of '8'
`define IN9 8'b00001001      // Encode of '9'
`define INA 8'b00001010      // Encode of 'A'
`define INB 8'b00001011      // Encode of 'B'
`define INC 8'b00001100      // Encode of 'C'
`define IND 8'b00001101      // Encode of 'D'
`define INE 8'b00001110      // Encode of 'E'
`define INF 8'b00001111      // Encode of 'F'
