module Forward (

);

endmodule