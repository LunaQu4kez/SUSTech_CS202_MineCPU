module BRU (
	input  logic [`DATA_WID] src1, src2,
	input  logic [`BRU_OP  ] op,
	output logic [`DATA_WID] res
);
	
endmodule