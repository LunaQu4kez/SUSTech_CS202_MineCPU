`include "Const.svh"

module ALU_Ctrl(
    input  [1:0] ALUop,
    input  [2:0] funct3,
    input  [6:0] funct7,
    output [3:0] ALUcontrol
);


endmodule