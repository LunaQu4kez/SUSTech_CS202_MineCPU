`include "Const.svh"

module Stage_WB (

);

endmodule