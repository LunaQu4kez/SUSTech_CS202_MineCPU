`include "Const.svh"

module Memory (
    
);




endmodule