`include "Const.svh"

module Stage_EX(

);
// TO-DO
	
endmodule