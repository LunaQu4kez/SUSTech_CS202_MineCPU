`define SEG_FREQ 200000                         // 500kHz
`define SEG0 8'b1111_1100                       // Display '0'
`define SEG1 8'b0110_0000                       // Display '1'
`define SEG2 8'b1101_1010                       // Display '2'
`define SEG3 8'b1111_0010                       // Display '3'
`define SEG4 8'b0110_0110                       // Display '4'
`define SEG5 8'b1011_0110                       // Display '5'
`define SEG6 8'b1011_1110                       // Display '6'
`define SEG7 8'b1110_0000                       // Display '7'
`define SEG8 8'b1111_1110                       // Display '8'
`define SEG9 8'b1111_0110                       // Display '9'
`define SEGA 8'b1110_1110                       // Display 'A'
`define SEGB 8'b0011_1110                       // Display 'B'
`define SEGC 8'b1001_1100                       // Display 'C'
`define SEGD 8'b0111_1010                       // Display 'D'
`define SEGE 8'b1001_1110                       // Display 'E'
`define SEGF 8'b1000_1110                       // Display 'F'
`define SEGH 8'b0110_1110                       // Display 'H'
`define SEGL 8'b0001_1100                       // Display 'L'
`define SEGo 8'b0011_1010                       // Display 'o'
`define SEGR 8'b0000_1010                       // Display 'r'
`define SEGt 8'b0001_1110                       // Display 't'
`define SEGu 8'b0011_1000                       // Display 'u'
`define SEGn 8'b0010_1010                       // Display 'n'
`define SEGN 8'b1110_1100                       // Display 'N'
`define SEGU 8'b0111_1100                       // Display 'U'
`define IN0 5'b00000                            // Encode of '0'
`define IN1 5'b00001                            // Encode of '1'
`define IN2 5'b00010                            // Encode of '2'
`define IN3 5'b00011                            // Encode of '3'
`define IN4 5'b00100                            // Encode of '4'
`define IN5 5'b00101                            // Encode of '5'
`define IN6 5'b00110                            // Encode of '6'
`define IN7 5'b00111                            // Encode of '7'
`define IN8 5'b01000                            // Encode of '8'
`define IN9 5'b01001                            // Encode of '9'
`define INA 5'b01010                            // Encode of 'A'
`define INB 5'b01011                            // Encode of 'B'
`define INC 5'b01100                            // Encode of 'C'
`define IND 5'b01101                            // Encode of 'D'
`define INE 5'b01110                            // Encode of 'E'
`define INF 5'b01111                            // Encode of 'F'
`define INH 5'b10000                            // Encode of 'H'
`define INL 5'b10001                            // Encode of 'L'
`define INo 5'b10010                            // Encode of 'o'
`define INR 5'b10011                            // Encode of 'r'
`define INt 5'b10100                            // Encode of 't'
`define INu 5'b10101                            // Encode of 'u'
`define INn 5'b10110                            // Encode of 'n'
`define INN 5'b10111                            // Encode of 'N'
`define INU 5'b11000                            // Encode of 'U'