`include "Const.svh"

module DCache (
    input logic             clk, rst,
);
    
endmodule
