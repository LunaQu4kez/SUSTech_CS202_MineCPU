`include "Const.svh"

module Stage_IF (

);

endmodule