`include "Const.svh"

module PC (
    input                    clk, rst,
    input  logic             PC_Write,   // hazard stall 1: yes, 0: no
    input  logic [`DATA_WID] new_pc,     // next pc
    output logic [`DATA_WID] pc_out
);

    logic [`DATA_WID] pc /*verilator public*/;
    assign pc_out = pc;

    initial pc = 0;

    always_ff @(negedge clk) begin
        if (rst) pc <= 0;
        else pc <= (PC_Write == 1'b0) ? new_pc : pc;
    end
    
endmodule
