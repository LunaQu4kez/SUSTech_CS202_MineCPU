`include "Const.svh"

module InstMem (
    input              clk,
    input  [`DATA_WID] addr,
    output [`DATA_WID] inst
);

    
    
endmodule
