`include "Const.svh"

module Stage_MEM (

);

endmodule